library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
 
entity rom is
generic(
    gADDRESS_WIDTH: natural := 12;
    gDATA_WIDTH: natural := 12
);
port(
    clock: in std_logic;
    rom_enable: in std_logic;
    address: in std_logic_vector((gADDRESS_WIDTH - 1) downto 0);
    data_output: out std_logic_vector ((gDATA_WIDTH - 1) downto 0)
);
end rom;
 
architecture arch of rom is
    --type rom_type is array (0 to (2**(gADDRESS_WIDTH) -1)) of std_logic_vector((gDATA_WIDTH - 1) downto 0);
    type rom_type is array (0 to (541 -1)) of std_logic_vector((gDATA_WIDTH - 1) downto 0);
    
    -- set the data on each adress to some value)
    constant mem: rom_type:=
    (
        "001100000010",
        "010000010100",
        "001110110100",
        "010000010101",
        "010111111111",
        "000000000000",
        "000000100000",
        "000000001110",
        "000000010101",
        "000000001100",
        "000000011000",
        "000000010110",
        "000000001110",
        "000000101011",
        "000000000000",
        "000000001011",
        "000000001010",
        "000000001101",
        "000000101011",
        "000000000000",
        "000000011010",
        "000000011110",
        "000000010010",
        "000000011101",
        "000000101011",
        "000000000000",
        "001000000010",
        "010000000100",
        "001000000011",
        "010000000101",
        "000100000000",
        "100000000100",
        "001000000000",
        "010000000100",
        "001000000001",
        "010000000101",
        "001000000100",
        "001100101011",
        "010100000000",
        "100011111111",
        "001000000011",
        "001100000001",
        "010001110000",
        "100000000011",
        "001100000001",
        "010000010100",
        "001100011010",
        "010000010101",
        "010111111111",
        "000000000000",
        "100011111110",
        "001100000010",
        "010000010000",
        "100000000000",
        "001111000110",
        "010000010000",
        "100000000001",
        "001100000001",
        "010000010000",
        "100000000010",
        "001100010100",
        "010000010000",
        "100000000011",
        "001100000001",
        "010000010100",
        "001100011010",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000001",
        "010000010000",
        "100000000000",
        "001101010111",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000100",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000101",
        "100000000110",
        "001100000001",
        "010000010000",
        "100000000000",
        "001101101011",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000111",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "100011111110",
        "001000000110",
        "010000000100",
        "001000000101",
        "010000000101",
        "000100000000",
        "100000000111",
        "001100101001",
        "010000010000",
        "100011111111",
        "010000110000",
        "100011111111",
        "001100101010",
        "010000010000",
        "100011111111",
        "001100000010",
        "010000010000",
        "100011111101",
        "001000000111",
        "010001110000",
        "100011111111",
        "001100000011",
        "010000010000",
        "100011111101",
        "001000000111",
        "010001110000",
        "100011111111",
        "001100000000",
        "010000010000",
        "100011111101",
        "001100000001",
        "010000010100",
        "001110001110",
        "010000010101",
        "000000000000",
        "010010000000",
        "001111111111",
        "010100000000",
        "001100000001",
        "010000010100",
        "001100110010",
        "010000010101",
        "001100011010",
        "010100000000",
        "001100000000",
        "010000010100",
        "001100000000",
        "010000010101",
        "001000000101",
        "001111111111",
        "010100000000",
        "001100000001",
        "010001110000",
        "100000000101",
        "001100000001",
        "010000010100",
        "001101101011",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000000",
        "010000010000",
        "100000000101",
        "001000000110",
        "001100000001",
        "010001110000",
        "100000000110",
        "001100000001",
        "010000010100",
        "001101101011",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000001",
        "010000010000",
        "100000000000",
        "001111000110",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000100",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000101",
        "100000000110",
        "001100000001",
        "010000010000",
        "100000000000",
        "001111011010",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000111",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "100000001011",
        "001000000101",
        "100000000111",
        "001000001011",
        "000000000000",
        "100011111110",
        "001100101000",
        "010000010000",
        "100011111111",
        "000000000000",
        "010010000000",
        "001100000001",
        "010000010100",
        "001111100100",
        "010000010101",
        "001111111111",
        "010100000000",
        "001100101011",
        "010100000000",
        "001100000001",
        "010000010100",
        "001100110010",
        "010000010101",
        "001100011010",
        "010100000000",
        "100011111111",
        "100000010001",
        "001100000001",
        "010000010100",
        "001111111010",
        "010000010101",
        "000000000000",
        "010010000000",
        "001111111111",
        "010100000000",
        "100011111111",
        "001100000010",
        "010000010100",
        "001100000011",
        "010000010101",
        "000000000000",
        "010010000000",
        "001111111111",
        "010100000000",
        "100011111111",
        "100000001001",
        "001100000010",
        "010000010100",
        "001100001101",
        "010000010101",
        "000000000000",
        "010010000000",
        "001111111111",
        "010100000000",
        "100011111111",
        "100000001010",
        "001100000010",
        "010000010000",
        "100000000000",
        "001100100100",
        "010000010000",
        "100000000001",
        "001100000000",
        "010000010000",
        "100000000010",
        "001100001001",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000110",
        "010000000100",
        "001000000111",
        "010000000101",
        "001000010001",
        "010000000011",
        "001000000101",
        "011000000000",
        "001100000000",
        "010000010000",
        "100011111101",
        "001100000000",
        "010000010100",
        "001100000000",
        "010000010101",
        "001000000111",
        "001111111111",
        "010100000000",
        "001100000001",
        "010001110000",
        "100000000111",
        "001100000001",
        "010000010100",
        "001111011111",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000000",
        "010000010000",
        "100000000111",
        "001000011011",
        "001100000001",
        "010001110000",
        "100000000110",
        "001100000001",
        "010000010100",
        "001111011111",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000010",
        "010000010000",
        "100000000000",
        "001101011110",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000100",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000101",
        "100000000110",
        "001100000010",
        "010000010000",
        "100000000000",
        "001101110010",
        "010000010000",
        "100000000001",
        "001101000000",
        "010000010000",
        "100000000010",
        "001100000111",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010100",
        "001101111000",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000110",
        "010000000100",
        "001000000101",
        "010000000101",
        "010111111111",
        "000000000000",
        "001100000000",
        "010000010000",
        "100000000101",
        "001000000010",
        "010000000100",
        "001000000011",
        "010000000101",
        "000100000000",
        "100000000100",
        "000000000000",
        "001100000000",
        "010000010000",
        "100011111101",
        "001100000010",
        "010000010100",
        "001110100011",
        "010000010101",
        "001000000100",
        "001100000000",
        "010100000000",
        "001100000001",
        "010000010000",
        "100011111101",
        "001000000100",
        "001100000001",
        "010001110000",
        "100000000100",
        "001100000000",
        "010000010000",
        "100011111101",
        "001100010000",
        "001000000101",
        "010001110000",
        "100000000101",
        "001000000100",
        "001100000000",
        "010100000000",
        "001100000010",
        "010000010100",
        "001110000010",
        "010000010101",
        "010111111111",
        "000000000000",
        "001000000010",
        "010000000100",
        "001000000011",
        "001100000001",
        "010001110000",
        "010000000101",
        "000100000000",
        "010000000001",
        "001000000101",
        "010001110000",
        "100000000101",
        "001000000000",
        "010000000100",
        "001000000001",
        "010000000101",
        "010111111111",
        "000000000000",
        "001100000001",
        "010000010000",
        "100000000010",
        "001100000110",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010000",
        "100000000000",
        "001111000110",
        "010000010000",
        "100000000001",
        "001100000001",
        "010000010100",
        "001100011010",
        "010000010101",
        "010111111111",
        "000000000000",
        "001100000000",
        "010000010000",
        "100011111101",
        "100011111110",
        "001101000000",
        "010000010000",
        "100000000100",
        "001100000001",
        "010000010000",
        "100000000101",
        "000000000000",
        "001100000010",
        "010000010100",
        "001111010001",
        "010000010101",
        "010010000000",
        "100000000110",
        "001111111111",
        "010100000000",
        "001000000100",
        "010000000100",
        "001000000101",
        "010000000101",
        "001000000110",
        "011000000000",
        "001000000101",
        "001100000001",
        "010001110000",
        "100000000101",
        "001000000110",
        "001100000010",
        "010000010100",
        "001111110001",
        "010000010101",
        "001100101011",
        "010100000000",
        "100011111111",
        "001100000010",
        "010000010100",
        "001111010001",
        "010000010101",
        "010111111111",
        "000000000000",
        "001101000000",
        "010000010100",
        "001100000001",
        "010000010101",
        "000100000000",
        "001100000001",
        "010000010100",
        "001101000101",
        "010000010101",
        "001100001101",
        "010100000000",
        "001100000001",
        "010000010100",
        "001110110100",
        "010000010101",
        "001100010110",
        "010100000000",
        "001100000010",
        "010000010100",
        "001101001100",
        "010000010101",
        "001100001110",
        "010100000000",
        "100011111110",
        "001100000001",
        "010000010000",
        "100000000010",
        "001100001111",
        "010000010000",
        "100000000011",
        "001100000010",
        "010000010000",
        "100000000000",
        "001111000110",
        "010000010000",
        "100000000001",
        "001100000001",
        "010000010100",
        "001100011010",
        "010000010101",
        "010111111111",
        "000011111111",
        "000000000000",
        "111100000000"        
    );
begin
 
process(clock) is
begin
    if(rising_edge(clock) and rom_enable = '1') then
        if conv_integer(unsigned(address))>540 then
            --Return zero as this is hoe long the program is
            data_output <= (others => '0');
        else
            --Return Valid ROM data.
            data_output <= mem(conv_integer(unsigned(address)));
        end if;
    end if;
end process;
 
end arch;